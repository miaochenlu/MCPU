`timescale 1ns / 1ps

`define LB   3'b001
`define LBU  3'b010
`define LH   3'b011
`define LHU  3'b100
`define LW   3'b101

`define SB  2'b01
`define SH  2'b10
`define SW  2'b11


`define MEM_INDEX_MSB 10
`define MEM_INDEX_LSB 4