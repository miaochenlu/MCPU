`timescale 1ns / 1ps

module LSQ (
    input clk,
    input rst,
    input rollback,

    input [ 3:0] LSQOp,
    input [31:0] MemAddr,
);

endmodule