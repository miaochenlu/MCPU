`timescale 1ns / 1ps

module HazardDetect(
    input ROB_full
    
);


endmodule